/*
 * Copyright (c) 2024 Will Park
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_uwasic_onboarding_WillPark (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  wire [7:0] en_reg_out_7_0;
  wire [7:0] en_reg_out_15_8;
  wire [7:0] en_reg_pwm_7_0;
  wire [7:0] en_reg_pwm_15_8;
  wire [7:0] pwm_duty_cycle;

  assign uio_oe = 8'hFF; // Set all IOs to output

  // Instantiate the PWM module
  pwm_peripheral pwm_peripheral_inst (
    .clk(clk),
    .rst_n(rst_n),
    .en_reg_out_7_0(en_reg_out_7_0),
    .en_reg_out_15_8(en_reg_out_15_8),
    .en_reg_pwm_7_0(en_reg_pwm_7_0),
    .en_reg_pwm_15_8(en_reg_pwm_15_8),
    .pwm_duty_cycle(pwm_duty_cycle),
    .out({uio_out, uo_out})
  );

  // List all unused inputs to prevent warnings
  wire _unused = &{ena, ui_in[7:3], uio_in, 1'b0};
  
  wire SCLK, COPI, nCS;
  assign SCLK = ui_in[0];
  assign COPI = ui_in[1];
  assign nCS = ui_in[2];

  // CDC Registers
  reg COPI_1;

  spi spi_inst (
    .rst_n(rst_n),
    .SCLK(SCLK),
    .COPI(COPI_1),
    .nCS(nCS),
    .data0(en_reg_out_7_0),
    .data1(en_reg_out_15_8),
    .data2(en_reg_pwm_7_0),
    .data3(en_reg_pwm_15_8),
    .data4(pwm_duty_cycle)
  );

  always @ (posedge clk) begin

    COPI_1 <= COPI;

  end

endmodule